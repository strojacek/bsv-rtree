module top ()

endmodule
